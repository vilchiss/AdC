library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity control_unit is
  port(
    clk: in std_logic
  );
end control_unit;

architecture arch of control_unit is

end architecture;
