library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity internal_registers is
  port(
    clk ; in std_logic
  );
end internal_registers;

architecture arch of internal_registers is

end architecture;
